#include "../../main.h"

// 开始自动生成静态结构
//	name	type	length	auth	value

@.	vlist	0	r	{
	help	string	0	r	_help_help
	format	string	0	r	_help_format
	
	// 导出
	_HELP_ROOT	-export	.
}

